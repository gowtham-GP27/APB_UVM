`define num_of_txns 1000
